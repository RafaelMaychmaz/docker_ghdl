library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

configuration b_config of b is
  for b_archi2
    --
  end for;
end configuration b_config;

